 module input_buffer(
    input logic 
 );
	
 
 
 endmodule