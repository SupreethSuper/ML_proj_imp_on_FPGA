`ifndef GLOBAL_DEFINES_VH
`define GLOBAL_DEFINES_VH
//==================GUARD RAILS==============

`define ADDR_WIDTH 32
`define DATA_WIDTH 32


//======NO CODE BEYOND THIS POINT==================
//=========END OF GUARD RAILS========================



`endif