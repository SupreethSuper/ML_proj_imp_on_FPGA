`ifndef GLOBAL_PARAMS_VH
`define GLOBAL_PARAMS_VH


//=========IMPORTS=================

`include "GLOBAL_DEFINES.vh"

//=============END OF IMPORTS=========

parameter ADDR_WIDTH = `ADDR_WIDTH;
parameter DATA_WIDTH = `DATA_WIDTH;




//=======================DO NOT CODE BEYOND THIS POINT==========
//======================END OF GUARD RAILS======================
`endif