 module input_buffer();
 
	
 
 
 endmodule